.title KiCad schematic
.include "models/C2012C0G2E102J085AA_p.mod"
.include "models/C2012X7R2A104K125AA_p.mod"
.include "models/C2012X7R2E103K125AA_p.mod"
.include "models/C3216X5R1H106M160AB_p.mod"
.include "models/MAX4080F.FAM"
XU1 /RSP VCC NC_01 0 /VOCM NC_02 NC_03 /RSN MAX4080F
R2 VCC /VOUT {Rsense}
R1 VCC /VOUT {Rsense}
R3 VCC /RSP 20
R4 /VOUT /RSN 20
XU5 /RSP /RSN C2012C0G2E102J085AA_p
I1 /VOUT 0 {ILOAD}
XU2 VCC 0 C3216X5R1H106M160AB_p
XU3 VCC 0 C2012X7R2A104K125AA_p
R5 /VOCM /CURRENT_FEEDBACK 100
XU4 /CURRENT_FEEDBACK 0 C2012X7R2E103K125AA_p
V1 VCC 0 {VIN}
.end
